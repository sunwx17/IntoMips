module cpu(
    );
endmodule
